class ahb_monitor extends uvm_monitor;

    ahb_config cfg;

    // Analysis port for individual beats
    uvm_analysis_port#(ahb_sequence_item) beat_ap;
    // Analysis port for completed burst transactions
    uvm_analysis_port#(ahb_burst_transaction) burst_ap;

    `uvm_component_utils(ahb_monitor)

    // Internal pipeline register for address phase
    protected ahb_sequence_item addr_phase_tr;
    protected bit addr_phase_valid = 0;

    // FSM for burst collection
    typedef enum {IDLE, IN_BURST} state_e;
    state_e state = IDLE;
    ahb_burst_transaction burst_tr;
    int beats_left;
    hburst_e active_burst_type;
    bit [31:0] start_addr;

    function new(string name = "ahb_monitor", uvm_component parent = null);
        super.new(name, parent);
        beat_ap = new("beat_ap", this);
        burst_ap = new("burst_ap", this);
    endfunction

    virtual task run_phase(uvm_phase phase);
        forever begin
            @(cfg.vif.monitor_cb);

            // -----------------------------------------------------------------
            // -- Data Phase Processing
            // -- Combine address (from last cycle) with data (from this cycle)
            // -----------------------------------------------------------------
            if (addr_phase_valid && cfg.vif.monitor_cb.HREADY) begin
                ahb_sequence_item complete_beat = addr_phase_tr;
                addr_phase_valid = 0; // Consume the address phase

                if (complete_beat.HWRITE) begin
                    complete_beat.HWDATA = cfg.vif.monitor_cb.HWDATA;
                end else begin
                    complete_beat.HRDATA = cfg.vif.monitor_cb.HRDATA;
                end
                
                process_complete_beat(complete_beat);
            end

            // -----------------------------------------------------------------
            // -- Address Phase Processing
            // -- Capture the start of a new transfer
            // -----------------------------------------------------------------
            if (cfg.vif.monitor_cb.HSELx && cfg.vif.monitor_cb.HTRANS inside {NONSEQ, SEQ}) begin
                if (addr_phase_valid) begin
                    `uvm_error("AHB_PROTOCOL_ERROR", "New transfer started before previous data phase completed (HREADY was low)")
                end
                addr_phase_tr = ahb_sequence_item::type_id::create("addr_phase_tr");
                addr_phase_tr.HADDR  = cfg.vif.monitor_cb.HADDR;
                addr_phase_tr.HWRITE = cfg.vif.monitor_cb.HWRITE;
                addr_phase_tr.HSIZE  = cfg.vif.monitor_cb.HSIZE;
                addr_phase_tr.HTRANS = cfg.vif.monitor_cb.HTRANS;
                addr_phase_tr.HWSTRB = cfg.vif.monitor_cb.HWSTRB;
                addr_phase_tr.HBURST = cfg.vif.monitor_cb.HBURST;
                addr_phase_tr.HPROT  = cfg.vif.monitor_cb.HPROT;
                addr_phase_valid = 1;
            end
        end
    endtask

    virtual protected task process_complete_beat(ahb_sequence_item beat);
        // Publish every complete beat
        beat_ap.write(beat);

        // Process the beat in the context of the burst FSM
        case (state)
            IDLE: begin
                if (beat.HTRANS == SEQ) begin
                    `uvm_error("AHB_PROTOCOL_ERROR", "SEQ transfer outside of a burst sequence")
                    return;
                end

                if (beat.HBURST == SINGLE) begin
                    ahb_burst_transaction single_beat_burst = new("single_beat_burst");
                    single_beat_burst.beats.push_back(beat);
                    burst_ap.write(single_beat_burst);
                end else begin // Start of a multi-beat burst
                    burst_tr = new("burst_tr");
                    burst_tr.beats.push_back(beat);
                    beats_left = get_burst_length(beat.HBURST) - 1;
                    active_burst_type = beat.HBURST;
                    start_addr = beat.HADDR;
                    state = IN_BURST;
                end
            end

            IN_BURST: begin
                if (beat.HTRANS != SEQ) begin
                    `uvm_error("AHB_PROTOCOL_ERROR", $sformatf("Burst started at %h of type %s terminated unexpectedly with HTRANS=%s", start_addr, active_burst_type.name(), beat.HTRANS.name()))
                    burst_ap.write(burst_tr); // Publish partial burst
                    state = IDLE;
                    // TODO: Re-process the current beat as a new transaction if it was NONSEQ
                    return;
                end
                if (beat.HBURST != active_burst_type) begin
                     `uvm_error("AHB_PROTOCOL_ERROR", $sformatf("HBURST changed mid-burst at address %h", beat.HADDR))
                end

                burst_tr.beats.push_back(beat);
                beats_left--;

                if (beats_left <= 0) {
                    burst_ap.write(burst_tr);
                    state = IDLE;
                end
            end
        endcase
    endtask

    function int get_burst_length(hburst_e burst);
        case(burst)
            SINGLE: return 1;
            INCR4, WRAP4: return 4;
            INCR8, WRAP8: return 8;
            INCR16, WRAP16: return 16;
            INCR: return -1; // Undefined length
            default: return 1;
        endcase
    endfunction

endclass
