package ahb_pkg;

    import uvm_pkg::*;

    `include "uvm_macros.svh"

    `include "ahb_types.svh"
    `include "ahb_config.svh"

    `include "ahb_sequence_item.svh"
    `include "ahb_burst_transaction.svh"
    `include "ahb_single_write_sequence.svh"
    `include "ahb_single_read_sequence.svh"
    `include "ahb_incr4_write_read_sequence.svh"
    `include "ahb_sequencer.svh"
    `include "ahb_driver.svh"
    `include "ahb_monitor.svh"
    `include "ahb_agent.svh"
    `include "ahb_env.svh"

endpackage